magic
tech sky130A
magscale 1 2
timestamp 1769127197
<< locali >>
rect 170 1960 479 2039
rect -96 0 96 151
rect 1056 0 1248 141
rect -200 -14 1400 0
rect -200 -194 294 -14
rect 474 -194 1400 -14
rect -200 -200 1400 -194
rect -96 -201 96 -200
<< viali >>
rect 294 -194 474 -14
<< metal1 >>
rect 672 3706 1143 3898
rect 160 108 224 3358
rect 951 3056 1143 3706
rect 673 2864 1143 3056
rect 951 1519 1143 2864
rect 668 1327 1143 1519
rect 951 702 1143 1327
rect 288 600 480 680
rect 673 510 1143 702
rect 288 -8 480 304
rect 672 40 864 120
rect 282 -14 486 -8
rect 282 -194 294 -14
rect 474 -194 486 -14
rect 282 -200 486 -194
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
<< labels >>
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBNS_5U
port 1 nsew signal bidirectional
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 2 nsew ground bidirectional
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBPS_20U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
